dual_port_bram.sv